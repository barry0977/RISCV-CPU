`include "const.v"

module ALU(
    
);
endmodule