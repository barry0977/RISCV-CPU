module InsFetch(

);
endmodule